module top_module ( input logic in, output logic out );
	assign out = in;
endmodule
