module add16 ( input [15:0] a, input [15:0] b, input cin, output [15:0] sum, output cout );
    // Module body
endmodule

module top_module (
    input [31:0] a,
    input [31:0] b,
    input sub,
    output [31:0] sum
);
    wire carry;
    wire [31:0] b_new;

    // (b ^ sub) = (~b) if sub=1
    assign b_new = b ^ {32{sub}};

    add16 adder1 (
        .a(a[15:0]),
        .b(b_new[15:0]),
        .cin(sub),
        .sum(sum[15:0]),
        .cout(carry)
    );
    add16 adder2 (
        .a(a[31:16]),
        .b(b_new[31:16]),
        .cin(carry),
        .sum(sum[31:16]),
        .cout()
    );
endmodule
